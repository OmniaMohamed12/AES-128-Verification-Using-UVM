package AES_Pack;
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    `include "AES_Sequence_Item.svh"
    `include "AES_Sequences.svh"
    `include "AES_Sequencer.svh"
    `include "AES_Driver.svh"
    `include "AES_Monitor.svh"
    `include "AES_Reference_Model.svh"
    `include "AES_Scoreboard.svh"
    `include "AES_Subscriber.svh"
    `include "AES_Agent.svh"
    `include "AES_Env.svh"
    `include "AES_Test.svh"
endpackage